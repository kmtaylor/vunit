-- This Source Code Form is subject to the terms of the Mozilla Public
-- License, v. 2.0. If a copy of the MPL was not distributed with this file,
-- You can obtain one at http://mozilla.org/MPL/2.0/.
--
-- Copyright (c) 2014-2022, Lars Asplund lars.anders.asplund@gmail.com

package body logger_pkg is

  procedure info(msg : string;
                 line_num : natural := 0;
                 file_name : string := "") is
  begin
    report(msg);
  end procedure;

end package body;
